/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    // Map some inputs to control signals
    wire load      = ui_in[7];
    wire [7:0] din = ui_in[7:0];

    // Counter instance
    wire [7:0] count_val;

    counter_8bit u_counter (
        .clk(clk),
        .rst_n(rst_n),
        .load(load),
        .en(ena),
        .data_in(count_val),
        .q(uo_out)
    );




  assign uo_out  = ui_in + uio_in;
  assign uio_out = 0;
  assign uio_oe  = 0;

  wire _unused = &{ena, clk, rst_n, 1'b0};


endmodule
